! Analisis de un hibrido 3 dB 180 disenyado
! para una frecuencia de 3 GHz.

DIM

  FREQ GHZ
  RES OH
  LNG mm
  TIME PS
  ANG DEG

VAR

  Wani  =  0.7733
  Wpue  =  1.497
  Radio  =  13.55
  ANGcorto  =  60
  LONGpue  =  13.83
  LONGlar  =  10.84
  LONGcor  =  2.59
  Inglete  =  0.01

CKT

! Aquí vendría algo del tipo:
! MSUB ER = erel H = hs T=espMet RHO = rMet RGH = rug

! Nombre Compo.   N1   N2    N3    Propiedades;  Donde Ni son los nodos a los
!                                                que el componente está aso-
!                                                ciado.


  MLIN_PUERTA1     1     2            W^Wpue     L^LONGpue
  MTEE             2     3    20      W1^Wpue    W2^Wani            W3^Wani
  MCURVE           3     4            W^Wani     ANG^ANGcorto       RAD^Radio
  MTEE             4     5     9      W1^Wani    W2^Wpue            W3^Wani
  MLIN             5     6            W^Wpue     L^LONGlar
  MBEND            6     7            W^Wpue     ANG = -30          M^Inglete
  MLIN_PUERTA2     7     8            W^Wpue     L^LONGcor
  MCURVE           9    10            W^Wani     ANG^ANGcorto       RAD^Radio
  MTEE            10    11    15      W1^Wani    W2^Wpue            W3^Wani
  MLIN            11    12            W^Wpue     L^LONGlar
  MBEND           12    13            W^Wpue     ANG = 30           M^Inglete
  MLIN_PUERTA3    13    14            W^Wpue     L^LONGcor
  MCURVE          15    16            W^Wani     ANG^ANGcorto       RAD^Radio
  MTEE            16    17    19      W1^Wani    W2^Wpue            W3^Wani
  MLIN_PUERTA4    17    18            W^Wpue     L^LNGpue
  MCURVE          19    20            W^Wani     ANG = 180          RAD^Radio

  DEF4P           2     8    14   18    Hibrido

! Ahora una red generada con el modelo de hibrido disponible
! en TouchStone

! HYBRID         21    22   23   24     L = 0     GIB = 0     PIB = 180

! DEF4P          21    22   23   24     Modelo

FREQ

  SWEEP 1 5 0.01

GRID

  GR1 -20 0 1
  GR1A -180 180 20

OUT

  Hibrido DB[S11] GR1
  Hibrido DB[S12] GR1
  Hibrido DB[S14] GR1
  Hibrido ANG[S12] GR1A
  Hibrido ANG[S14] GR1A
  Hibrido s11 sc1
